library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	7846	)	,
(	7831	)	,
(	7815	)	,
(	7800	)	,
(	7784	)	,
(	7768	)	,
(	7753	)	,
(	7737	)	,
(	7722	)	,
(	7707	)	,
(	7691	)	,
(	7676	)	,
(	7660	)	,
(	7645	)	,
(	7630	)	,
(	7614	)	,
(	7599	)	,
(	7584	)	,
(	7569	)	,
(	7554	)	,
(	7538	)	,
(	7523	)	,
(	7508	)	,
(	7493	)	,
(	7478	)	,
(	7463	)	,
(	7448	)	,
(	7433	)	,
(	7418	)	,
(	7403	)	,
(	7388	)	,
(	7374	)	,
(	7359	)	,
(	7344	)	,
(	7329	)	,
(	7314	)	,
(	7300	)	,
(	7285	)	,
(	7270	)	,
(	7256	)	,
(	7241	)	,
(	7226	)	,
(	7212	)	,
(	7197	)	,
(	7183	)	,
(	7168	)	,
(	7154	)	,
(	7139	)	,
(	7125	)	,
(	7111	)	,
(	7096	)	,
(	7082	)	,
(	7067	)	,
(	7053	)	,
(	7039	)	,
(	7025	)	,
(	7010	)	,
(	6996	)	,
(	6982	)	,
(	6968	)	,
(	6954	)	,
(	6940	)	,
(	6926	)	,
(	6912	)	,
(	6898	)	,
(	6884	)	,
(	6870	)	,
(	6856	)	,
(	6842	)	,
(	6828	)	,
(	6814	)	,
(	6800	)	,
(	6787	)	,
(	6773	)	,
(	6759	)	,
(	6745	)	,
(	6732	)	,
(	6718	)	,
(	6704	)	,
(	6691	)	,
(	6677	)	,
(	6663	)	,
(	6650	)	,
(	6636	)	,
(	6623	)	,
(	6609	)	,
(	6596	)	,
(	6582	)	,
(	6569	)	,
(	6556	)	,
(	6542	)	,
(	6529	)	,
(	6516	)	,
(	6502	)	,
(	6489	)	,
(	6476	)	,
(	6463	)	,
(	6449	)	,
(	6436	)	,
(	6423	)	,
(	6410	)	,
(	6397	)	,
(	6384	)	,
(	6371	)	,
(	6358	)	,
(	6345	)	,
(	6332	)	,
(	6319	)	,
(	6306	)	,
(	6293	)	,
(	6280	)	,
(	6267	)	,
(	6254	)	,
(	6241	)	,
(	6229	)	,
(	6216	)	,
(	6203	)	,
(	6190	)	,
(	6178	)	,
(	6165	)	,
(	6152	)	,
(	6140	)	,
(	6127	)	,
(	6115	)	,
(	6102	)	,
(	6090	)	,
(	6077	)	,
(	6065	)	,
(	6052	)	,
(	6040	)	,
(	6027	)	,
(	6015	)	,
(	6003	)	,
(	5990	)	,
(	5978	)	,
(	5966	)	,
(	5953	)	,
(	5941	)	,
(	5929	)	,
(	5917	)	,
(	5905	)	,
(	5892	)	,
(	5880	)	,
(	5868	)	,
(	5856	)	,
(	5844	)	,
(	5832	)	,
(	5820	)	,
(	5808	)	,
(	5796	)	,
(	5784	)	,
(	5772	)	,
(	5760	)	,
(	5748	)	,
(	5736	)	,
(	5725	)	,
(	5713	)	,
(	5701	)	,
(	5689	)	,
(	5677	)	,
(	5666	)	,
(	5654	)	,
(	5642	)	,
(	5631	)	,
(	5619	)	,
(	5607	)	,
(	5596	)	,
(	5584	)	,
(	5573	)	,
(	5561	)	,
(	5550	)	,
(	5538	)	,
(	5527	)	,
(	5515	)	,
(	5504	)	,
(	5492	)	,
(	5481	)	,
(	5470	)	,
(	5458	)	,
(	5447	)	,
(	5436	)	,
(	5425	)	,
(	5413	)	,
(	5402	)	,
(	5391	)	,
(	5380	)	,
(	5369	)	,
(	5357	)	,
(	5346	)	,
(	5335	)	,
(	5324	)	,
(	5313	)	,
(	5302	)	,
(	5291	)	,
(	5280	)	,
(	5269	)	,
(	5258	)	,
(	5247	)	,
(	5236	)	,
(	5226	)	,
(	5215	)	,
(	5204	)	,
(	5193	)	,
(	5182	)	,
(	5172	)	,
(	5161	)	,
(	5150	)	,
(	5139	)	,
(	5129	)	,
(	5118	)	,
(	5107	)	,
(	5097	)	,
(	5086	)	,
(	5076	)	,
(	5065	)	,
(	5054	)	,
(	5044	)	,
(	5033	)	,
(	5023	)	,
(	5013	)	,
(	5002	)	,
(	4992	)	,
(	4981	)	,
(	4971	)	,
(	4961	)	,
(	4950	)	,
(	4940	)	,
(	4930	)	,
(	4919	)	,
(	4909	)	,
(	4899	)	,
(	4889	)	,
(	4879	)	,
(	4868	)	,
(	4858	)	,
(	4848	)	,
(	4838	)	,
(	4828	)	,
(	4818	)	,
(	4808	)	,
(	4798	)	,
(	4788	)	,
(	4778	)	,
(	4768	)	,
(	4758	)	,
(	4748	)	,
(	4738	)	,
(	4728	)	,
(	4718	)	,
(	4708	)	,
(	4699	)	,
(	4689	)	,
(	4679	)	,
(	4669	)	,
(	4660	)	,
(	4650	)	,
(	4640	)	,
(	4630	)	,
(	4621	)	,
(	4611	)	,
(	4601	)	,
(	4592	)	,
(	4582	)	,
(	4573	)	,
(	4563	)	,
(	4554	)	,
(	4544	)	,
(	4535	)	,
(	4525	)	,
(	4516	)	,
(	4506	)	,
(	4497	)	,
(	4487	)	,
(	4478	)	,
(	4469	)	,
(	4459	)	,
(	4450	)	,
(	4441	)	,
(	4432	)	,
(	4422	)	,
(	4413	)	,
(	4404	)	,
(	4395	)	,
(	4385	)	,
(	4376	)	,
(	4367	)	,
(	4358	)	,
(	4349	)	,
(	4340	)	,
(	4331	)	,
(	4322	)	,
(	4313	)	,
(	4304	)	,
(	4295	)	,
(	4286	)	,
(	4277	)	,
(	4268	)	,
(	4259	)	,
(	4250	)	,
(	4241	)	,
(	4232	)	,
(	4223	)	,
(	4215	)	,
(	4206	)	,
(	4197	)	,
(	4188	)	,
(	4179	)	,
(	4171	)	,
(	4162	)	,
(	4153	)	,
(	4145	)	,
(	4136	)	,
(	4127	)	,
(	4119	)	,
(	4110	)	,
(	4101	)	,
(	4093	)	,
(	4084	)	,
(	4076	)	,
(	4067	)	,
(	4059	)	,
(	4050	)	,
(	4042	)	,
(	4033	)	,
(	4025	)	,
(	4017	)	,
(	4008	)	,
(	4000	)	,
(	3991	)	,
(	3983	)	,
(	3975	)	,
(	3967	)	,
(	3958	)	,
(	3950	)	,
(	3942	)	,
(	3933	)	,
(	3925	)	,
(	3917	)	,
(	3909	)	,
(	3901	)	,
(	3893	)	,
(	3884	)	,
(	3876	)	,
(	3868	)	,
(	3860	)	,
(	3852	)	,
(	3844	)	,
(	3836	)	,
(	3828	)	,
(	3820	)	,
(	3812	)	,
(	3804	)	,
(	3796	)	,
(	3788	)	,
(	3780	)	,
(	3773	)	,
(	3765	)	,
(	3757	)	,
(	3749	)	,
(	3741	)	,
(	3733	)	,
(	3726	)	,
(	3718	)	,
(	3710	)	,
(	3702	)	,
(	3695	)	,
(	3687	)	,
(	3679	)	,
(	3672	)	,
(	3664	)	,
(	3656	)	,
(	3649	)	,
(	3641	)	,
(	3634	)	,
(	3626	)	,
(	3619	)	,
(	3611	)	,
(	3603	)	,
(	3596	)	,
(	3589	)	,
(	3581	)	,
(	3574	)	,
(	3566	)	,
(	3559	)	,
(	3551	)	,
(	3544	)	,
(	3537	)	,
(	3529	)	,
(	3522	)	,
(	3515	)	,
(	3507	)	,
(	3500	)	,
(	3493	)	,
(	3486	)	,
(	3478	)	,
(	3471	)	,
(	3464	)	,
(	3457	)	,
(	3450	)	,
(	3442	)	,
(	3435	)	,
(	3428	)	,
(	3421	)	,
(	3414	)	,
(	3407	)	,
(	3400	)	,
(	3393	)	,
(	3386	)	,
(	3379	)	,
(	3372	)	,
(	3365	)	,
(	3358	)	,
(	3351	)	,
(	3344	)	,
(	3337	)	,
(	3330	)	,
(	3323	)	,
(	3316	)	,
(	3310	)	,
(	3303	)	,
(	3296	)	,
(	3289	)	,
(	3282	)	,
(	3276	)	,
(	3269	)	,
(	3262	)	,
(	3255	)	,
(	3249	)	,
(	3242	)	,
(	3235	)	,
(	3229	)	,
(	3222	)	,
(	3215	)	,
(	3209	)	,
(	3202	)	,
(	3195	)	,
(	3189	)	,
(	3182	)	,
(	3176	)	,
(	3169	)	,
(	3163	)	,
(	3156	)	,
(	3150	)	,
(	3143	)	,
(	3137	)	,
(	3130	)	,
(	3124	)	,
(	3118	)	,
(	3111	)	,
(	3105	)	,
(	3098	)	,
(	3092	)	,
(	3086	)	,
(	3079	)	,
(	3073	)	,
(	3067	)	,
(	3061	)	,
(	3054	)	,
(	3048	)	,
(	3042	)	,
(	3036	)	,
(	3029	)	,
(	3023	)	,
(	3017	)	,
(	3011	)	,
(	3005	)	,
(	2999	)	,
(	2993	)	,
(	2986	)	,
(	2980	)	,
(	2974	)	,
(	2968	)	,
(	2962	)	,
(	2956	)	,
(	2950	)	,
(	2944	)	,
(	2938	)	,
(	2932	)	,
(	2926	)	,
(	2920	)	,
(	2914	)	,
(	2908	)	,
(	2902	)	,
(	2897	)	,
(	2891	)	,
(	2885	)	,
(	2879	)	,
(	2873	)	,
(	2867	)	,
(	2862	)	,
(	2856	)	,
(	2850	)	,
(	2844	)	,
(	2839	)	,
(	2833	)	,
(	2827	)	,
(	2821	)	,
(	2816	)	,
(	2810	)	,
(	2804	)	,
(	2799	)	,
(	2793	)	,
(	2787	)	,
(	2782	)	,
(	2776	)	,
(	2771	)	,
(	2765	)	,
(	2759	)	,
(	2754	)	,
(	2748	)	,
(	2743	)	,
(	2737	)	,
(	2732	)	,
(	2726	)	,
(	2721	)	,
(	2716	)	,
(	2710	)	,
(	2705	)	,
(	2699	)	,
(	2694	)	,
(	2688	)	,
(	2683	)	,
(	2678	)	,
(	2672	)	,
(	2667	)	,
(	2662	)	,
(	2656	)	,
(	2651	)	,
(	2646	)	,
(	2641	)	,
(	2635	)	,
(	2630	)	,
(	2625	)	,
(	2620	)	,
(	2614	)	,
(	2609	)	,
(	2604	)	,
(	2599	)	,
(	2594	)	,
(	2589	)	,
(	2584	)	,
(	2578	)	,
(	2573	)	,
(	2568	)	,
(	2563	)	,
(	2558	)	,
(	2553	)	,
(	2548	)	,
(	2543	)	,
(	2538	)	,
(	2533	)	,
(	2528	)	,
(	2523	)	,
(	2518	)	,
(	2513	)	,
(	2508	)	,
(	2503	)	,
(	2498	)	,
(	2494	)	,
(	2489	)	,
(	2484	)	,
(	2479	)	,
(	2474	)	,
(	2469	)	,
(	2464	)	,
(	2460	)	,
(	2455	)	,
(	2450	)	,
(	2445	)	,
(	2440	)	,
(	2436	)	,
(	2431	)	,
(	2426	)	,
(	2422	)	,
(	2417	)	,
(	2412	)	,
(	2408	)	,
(	2403	)	,
(	2398	)	,
(	2394	)	,
(	2389	)	,
(	2384	)	,
(	2380	)	,
(	2375	)	,
(	2371	)	,
(	2366	)	,
(	2361	)	,
(	2357	)	,
(	2352	)	,
(	2348	)	,
(	2343	)	,
(	2339	)	,
(	2334	)	,
(	2330	)	,
(	2325	)	,
(	2321	)	,
(	2316	)	,
(	2312	)	,
(	2308	)	,
(	2303	)	,
(	2299	)	,
(	2294	)	,
(	2290	)	,
(	2286	)	,
(	2281	)	,
(	2277	)	,
(	2273	)	,
(	2268	)	,
(	2264	)	,
(	2260	)	,
(	2256	)	,
(	2251	)	,
(	2247	)	,
(	2243	)	,
(	2238	)	,
(	2234	)	,
(	2230	)	,
(	2226	)	,
(	2222	)	,
(	2217	)	,
(	2213	)	,
(	2209	)	,
(	2205	)	,
(	2201	)	,
(	2197	)	,
(	2193	)	,
(	2189	)	,
(	2184	)	,
(	2180	)	,
(	2176	)	,
(	2172	)	,
(	2168	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2152	)	,
(	2148	)	,
(	2144	)	,
(	2140	)	,
(	2136	)	,
(	2132	)	,
(	2128	)	,
(	2124	)	,
(	2120	)	,
(	2117	)	,
(	2113	)	,
(	2109	)	,
(	2105	)	,
(	2101	)	,
(	2097	)	,
(	2093	)	,
(	2089	)	,
(	2086	)	,
(	2082	)	,
(	2078	)	,
(	2074	)	,
(	2070	)	,
(	2067	)	,
(	2063	)	,
(	2059	)	,
(	2055	)	,
(	2052	)	,
(	2048	)	,
(	2044	)	,
(	2041	)	,
(	2037	)	,
(	2033	)	,
(	2030	)	,
(	2026	)	,
(	2022	)	,
(	2019	)	,
(	2015	)	,
(	2011	)	,
(	2008	)	,
(	2004	)	,
(	2001	)	,
(	1997	)	,
(	1993	)	,
(	1990	)	,
(	1986	)	,
(	1983	)	,
(	1979	)	,
(	1976	)	,
(	1972	)	,
(	1969	)	,
(	1965	)	,
(	1962	)	,
(	1958	)	,
(	1955	)	,
(	1951	)	,
(	1948	)	,
(	1944	)	,
(	1941	)	,
(	1938	)	,
(	1934	)	,
(	1931	)	,
(	1927	)	,
(	1924	)	,
(	1921	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1907	)	,
(	1904	)	,
(	1901	)	,
(	1897	)	,
(	1894	)	,
(	1891	)	,
(	1888	)	,
(	1884	)	,
(	1881	)	,
(	1878	)	,
(	1875	)	,
(	1871	)	,
(	1868	)	,
(	1865	)	,
(	1862	)	,
(	1858	)	,
(	1855	)	,
(	1852	)	,
(	1849	)	,
(	1846	)	,
(	1843	)	,
(	1840	)	,
(	1836	)	,
(	1833	)	,
(	1830	)	,
(	1827	)	,
(	1824	)	,
(	1821	)	,
(	1818	)	,
(	1815	)	,
(	1812	)	,
(	1809	)	,
(	1806	)	,
(	1803	)	,
(	1800	)	,
(	1797	)	,
(	1794	)	,
(	1791	)	,
(	1788	)	,
(	1785	)	,
(	1782	)	,
(	1779	)	,
(	1776	)	,
(	1773	)	,
(	1770	)	,
(	1767	)	,
(	1764	)	,
(	1761	)	,
(	1758	)	,
(	1755	)	,
(	1753	)	,
(	1750	)	,
(	1747	)	,
(	1744	)	,
(	1741	)	,
(	1738	)	,
(	1735	)	,
(	1733	)	,
(	1730	)	,
(	1727	)	,
(	1724	)	,
(	1721	)	,
(	1719	)	,
(	1716	)	,
(	1713	)	,
(	1710	)	,
(	1708	)	,
(	1705	)	,
(	1702	)	,
(	1699	)	,
(	1697	)	,
(	1694	)	,
(	1691	)	,
(	1689	)	,
(	1686	)	,
(	1683	)	,
(	1681	)	,
(	1678	)	,
(	1675	)	,
(	1673	)	,
(	1670	)	,
(	1667	)	,
(	1665	)	,
(	1662	)	,
(	1660	)	,
(	1657	)	,
(	1654	)	,
(	1652	)	,
(	1649	)	,
(	1647	)	,
(	1644	)	,
(	1642	)	,
(	1639	)	,
(	1637	)	,
(	1634	)	,
(	1632	)	,
(	1629	)	,
(	1627	)	,
(	1624	)	,
(	1622	)	,
(	1619	)	,
(	1617	)	,
(	1614	)	,
(	1612	)	,
(	1609	)	,
(	1607	)	,
(	1604	)	,
(	1602	)	,
(	1600	)	,
(	1597	)	,
(	1595	)	,
(	1592	)	,
(	1590	)	,
(	1588	)	,
(	1585	)	,
(	1583	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1573	)	,
(	1571	)	,
(	1569	)	,
(	1567	)	,
(	1564	)	,
(	1562	)	,
(	1560	)	,
(	1557	)	,
(	1555	)	,
(	1553	)	,
(	1551	)	,
(	1548	)	,
(	1546	)	,
(	1544	)	,
(	1542	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1533	)	,
(	1530	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1517	)	,
(	1515	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1507	)	,
(	1505	)	,
(	1503	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1494	)	,
(	1492	)	,
(	1490	)	,
(	1488	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1480	)	,
(	1478	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1460	)	,
(	1458	)	,
(	1456	)	,
(	1454	)	,
(	1452	)	,
(	1450	)	,
(	1448	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1440	)	,
(	1439	)	,
(	1437	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1427	)	,
(	1425	)	,
(	1424	)	,
(	1422	)	,
(	1420	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1407	)	,
(	1405	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1398	)	,
(	1397	)	,
(	1395	)	,
(	1393	)	,
(	1391	)	,
(	1390	)	,
(	1388	)	,
(	1386	)	,
(	1384	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1378	)	,
(	1376	)	,
(	1374	)	,
(	1372	)	,
(	1371	)	,
(	1369	)	,
(	1367	)	,
(	1366	)	,
(	1364	)	,
(	1362	)	,
(	1361	)	,
(	1359	)	,
(	1358	)	,
(	1356	)	,
(	1354	)	,
(	1353	)	,
(	1351	)	,
(	1350	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1338	)	,
(	1337	)	,
(	1335	)	,
(	1334	)	,
(	1332	)	,
(	1331	)	,
(	1329	)	,
(	1328	)	,
(	1326	)	,
(	1325	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1319	)	,
(	1317	)	,
(	1316	)	,
(	1314	)	,
(	1313	)	,
(	1311	)	,
(	1310	)	,
(	1308	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1295	)	,
(	1294	)	,
(	1293	)	,
(	1291	)	,
(	1290	)	,
(	1288	)	,
(	1287	)	,
(	1286	)	,
(	1284	)	,
(	1283	)	,
(	1281	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1272	)	,
(	1271	)	,
(	1269	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1253	)	,
(	1251	)	,
(	1250	)	,
(	1249	)	,
(	1248	)	,
(	1246	)	,
(	1245	)	,
(	1244	)	,
(	1243	)	,
(	1241	)	,
(	1240	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1235	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1230	)	,
(	1229	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1220	)	,
(	1219	)	,
(	1218	)	,
(	1217	)	,
(	1215	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1208	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1166	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1157	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1077	)	,
(	1076	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1070	)	,
(	1069	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1067	)	,
(	1066	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1064	)	,
(	1063	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1061	)	,
(	1060	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1058	)	,
(	1057	)	,
(	1057	)	,
(	1056	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1054	)	,
(	1053	)	,
(	1053	)	,
(	1052	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1050	)	,
(	1049	)	,
(	1049	)	,
(	1048	)	,
(	1048	)	,
(	1047	)	,
(	1047	)	,
(	1046	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1044	)	,
(	1043	)	,
(	1043	)	,
(	1042	)	,
(	1042	)	,
(	1041	)	,
(	1041	)	,
(	1040	)	,
(	1040	)	,
(	1039	)	,
(	1039	)	,
(	1038	)	,
(	1038	)	,
(	1037	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1035	)	,
(	1034	)	,
(	1034	)	,
(	1033	)	,
(	1033	)	,
(	1032	)	,
(	1032	)	,
(	1031	)	,
(	1031	)	,
(	1030	)	,
(	1030	)	,
(	1029	)	,
(	1029	)	,
(	1028	)	,
(	1028	)	,
(	1027	)	,
(	1027	)	,
(	1026	)	,
(	1026	)	,
(	1025	)	,
(	1025	)	,
(	1025	)	,
(	1024	)	,
(	1024	)	,
(	1023	)	,
(	1023	)	,
(	1022	)	,
(	1022	)	,
(	1021	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1019	)	,
(	1018	)	,
(	1018	)	,
(	1017	)	,
(	1017	)	,
(	1016	)	,
(	1016	)	,
(	1015	)	,
(	1015	)	,
(	1015	)	,
(	1014	)	,
(	1014	)	,
(	1013	)	,
(	1013	)	,
(	1012	)	,
(	1012	)	,
(	1011	)	,
(	1011	)	,
(	1010	)	,
(	1010	)	,
(	1010	)	,
(	1009	)	,
(	1009	)	,
(	1008	)	,
(	1008	)	,
(	1007	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1005	)	,
(	1004	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1002	)	,
(	1002	)	,
(	1001	)	,
(	1001	)	,
(	1000	)	,
(	1000	)	,
(	999	)	,
(	999	)	,
(	999	)	,
(	998	)	,
(	998	)	,
(	997	)	,
(	997	)	,
(	996	)	,
(	996	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	994	)	,
(	993	)	,
(	993	)	,
(	993	)	,
(	992	)	,
(	992	)	,
(	991	)	,
(	991	)	,
(	991	)	,
(	990	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	988	)	,
(	988	)	,
(	987	)	,
(	987	)	,
(	986	)	,
(	986	)	,
(	986	)	,
(	985	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	983	)	,
(	982	)	,
(	982	)	,
(	981	)	,
(	981	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	979	)	,
(	979	)	,
(	978	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	974	)	,
(	973	)	,
(	973	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	971	)	,
(	971	)	,
(	970	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	966	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	964	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	953	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	951	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	949	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	947	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	940	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	934	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	666	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	612	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	576	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	554	)	,
(	553	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	543	)	,
(	542	)	,
(	541	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	513	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	509	)	,
(	508	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	503	)	,
(	502	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	498	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	492	)	,
(	491	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	487	)	,
(	486	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	482	)	,
(	481	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	477	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	472	)	,
(	471	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	467	)	,
(	466	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	462	)	,
(	461	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	457	)	,
(	456	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	452	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	448	)	,
(	447	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	443	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	439	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	435	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	431	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	427	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	423	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	419	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	412	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	405	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	362	)	,
(	361	)	,
(	361	)	,
(	360	)	,
(	359	)	,
(	359	)	,
(	358	)	,
(	357	)	,
(	357	)	,
(	356	)	,
(	355	)	,
(	355	)	,
(	354	)	,
(	353	)	,
(	353	)	,
(	352	)	,
(	351	)	,
(	351	)	,
(	350	)	,
(	349	)	,
(	349	)	,
(	348	)	,
(	347	)	,
(	347	)	,
(	346	)	,
(	345	)	,
(	345	)	,
(	344	)	,
(	343	)	,
(	343	)	,
(	342	)	,
(	342	)	,
(	341	)	,
(	340	)	,
(	340	)	,
(	339	)	,
(	338	)	,
(	338	)	,
(	337	)	,
(	337	)	,
(	336	)	,
(	335	)	,
(	335	)	,
(	334	)	,
(	334	)	,
(	333	)	,
(	332	)	,
(	332	)	,
(	331	)	,
(	331	)	,
(	330	)	,
(	329	)	,
(	329	)	,
(	328	)	,
(	328	)	,
(	327	)	,
(	326	)	,
(	326	)	,
(	325	)	,
(	325	)	,
(	324	)	,
(	324	)	,
(	323	)	,
(	322	)	,
(	322	)	,
(	321	)	,
(	321	)	,
(	320	)	,
(	320	)	,
(	319	)	,
(	319	)	,
(	318	)	,
(	318	)	,
(	317	)	,
(	316	)	,
(	316	)	,
(	315	)	,
(	315	)	,
(	314	)	,
(	314	)	,
(	313	)	,
(	313	)	,
(	312	)	,
(	312	)	,
(	311	)	,
(	311	)	,
(	310	)	,
(	310	)	,
(	309	)	,
(	309	)	,
(	308	)	,
(	308	)	,
(	307	)	,
(	307	)	,
(	306	)	,
(	306	)	,
(	305	)	,
(	305	)	,
(	304	)	,
(	304	)	,
(	303	)	,
(	303	)	,
(	303	)	,
(	302	)	,
(	302	)	,
(	301	)	,
(	301	)	,
(	300	)	,
(	300	)	,
(	299	)	,
(	299	)	,
(	298	)	,
(	298	)	,
(	298	)	,
(	297	)	,
(	297	)	,
(	296	)	,
(	296	)	,
(	296	)	,
(	295	)	,
(	295	)	,
(	294	)	,
(	294	)	,
(	293	)	,
(	293	)	,
(	293	)	,
(	292	)	,
(	292	)	,
(	291	)	,
(	291	)	,
(	291	)	,
(	290	)	,
(	290	)	,
(	290	)	,
(	289	)	,
(	289	)	,
(	289	)	,
(	288	)	,
(	288	)	,
(	287	)	,
(	287	)	,
(	287	)	,
(	286	)	,
(	286	)	,
(	286	)	,
(	285	)	,
(	285	)	,
(	285	)	,
(	284	)	,
(	284	)	,
(	284	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	282	)	,
(	282	)	,
(	282	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	280	)	,
(	280	)	,
(	280	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	270	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	271	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	272	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	273	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	274	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	275	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	276	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	277	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	278	)	,
(	279	)	,
(	279	)	,
(	279	)	,
(	280	)	,
(	280	)	,
(	280	)	,
(	280	)	,
(	281	)	,
(	281	)	,
(	281	)	,
(	282	)	,
(	282	)	,
(	283	)	,
(	283	)	,
(	283	)	,
(	284	)	,
(	284	)	,
(	284	)	,
(	285	)	,
(	285	)	,
(	286	)	,
(	286	)	,
(	286	)	,
(	287	)	,
(	287	)	,
(	288	)	,
(	288	)	,
(	288	)	,
(	289	)	,
(	289	)	,
(	290	)	,
(	290	)	,
(	291	)	,
(	291	)	,
(	292	)	,
(	292	)	,
(	293	)	,
(	293	)	,
(	294	)	,
(	294	)	,
(	295	)	,
(	295	)	,
(	296	)	,
(	296	)	,
(	297	)	,
(	297	)	,
(	298	)	,
(	298	)	,
(	299	)	,
(	299	)	,
(	300	)	,
(	301	)	,
(	301	)	,
(	302	)	,
(	302	)	,
(	303	)	,
(	304	)	,
(	304	)	,
(	305	)	,
(	305	)	,
(	306	)	,
(	307	)	,
(	307	)	,
(	308	)	,
(	309	)	,
(	309	)	,
(	310	)	,
(	311	)	,
(	311	)	,
(	312	)	,
(	313	)	,
(	313	)	,
(	314	)	,
(	315	)	,
(	315	)	,
(	316	)	,
(	317	)	,
(	318	)	,
(	318	)	,
(	319	)	,
(	320	)	,
(	321	)	,
(	321	)	,
(	322	)	,
(	323	)	,
(	324	)	,
(	325	)	,
(	325	)	,
(	326	)	,
(	327	)	,
(	328	)	,
(	329	)	,
(	329	)	,
(	330	)	,
(	331	)	,
(	332	)	,
(	333	)	,
(	334	)	,
(	335	)	,
(	336	)	,
(	336	)	,
(	337	)	,
(	338	)	,
(	339	)	,
(	340	)	,
(	341	)	,
(	342	)	,
(	343	)	,
(	344	)	,
(	345	)	,
(	346	)	,
(	347	)	,
(	348	)	,
(	349	)	,
(	350	)	,
(	351	)	,
(	352	)	,
(	353	)	,
(	354	)	,
(	355	)	,
(	356	)	,
(	357	)	,
(	358	)	,
(	359	)	,
(	360	)	,
(	361	)	,
(	362	)	,
(	363	)	,
(	364	)	,
(	365	)	,
(	366	)	,
(	367	)	,
(	369	)	,
(	370	)	,
(	371	)	,
(	372	)	,
(	373	)	,
(	374	)	,
(	375	)	,
(	377	)	,
(	378	)	,
(	379	)	,
(	380	)	,
(	381	)	,
(	382	)	,
(	384	)	,
(	385	)	,
(	386	)	,
(	387	)	,
(	389	)	,
(	390	)	,
(	391	)	,
(	392	)	,
(	394	)	,
(	395	)	,
(	396	)	,
(	398	)	,
(	399	)	,
(	400	)	,
(	401	)	,
(	403	)	,
(	404	)	,
(	405	)	,
(	407	)	,
(	408	)	,
(	410	)	,
(	411	)	,
(	412	)	,
(	414	)	,
(	415	)	,
(	416	)	,
(	418	)	,
(	419	)	,
(	421	)	,
(	422	)	,
(	424	)	,
(	425	)	,
(	427	)	,
(	428	)	,
(	429	)	,
(	431	)	,
(	432	)	,
(	434	)	,
(	435	)	,
(	437	)	,
(	439	)	,
(	440	)	,
(	442	)	,
(	443	)	,
(	445	)	,
(	446	)	,
(	448	)	,
(	449	)	,
(	451	)	,
(	453	)	,
(	454	)	,
(	456	)	,
(	458	)	,
(	459	)	,
(	461	)	,
(	462	)	,
(	464	)	,
(	466	)	,
(	467	)	,
(	469	)	,
(	471	)	,
(	473	)	,
(	474	)	,
(	476	)	,
(	478	)	,
(	479	)	,
(	481	)	,
(	483	)	,
(	485	)	,
(	487	)	,
(	488	)	,
(	490	)	,
(	492	)	,
(	494	)	,
(	496	)	,
(	497	)	,
(	499	)	,
(	501	)	,
(	503	)	,
(	505	)	,
(	507	)	,
(	509	)	,
(	510	)	,
(	512	)	,
(	514	)	,
(	516	)	,
(	518	)	,
(	520	)	,
(	522	)	,
(	524	)	,
(	526	)	,
(	528	)	,
(	530	)	,
(	532	)	,
(	534	)	,
(	536	)	,
(	538	)	,
(	540	)	,
(	542	)	,
(	544	)	,
(	546	)	,
(	548	)	,
(	550	)	,
(	552	)	,
(	554	)	,
(	557	)	,
(	559	)	,
(	561	)	,
(	563	)	,
(	565	)	,
(	567	)	,
(	569	)	,
(	572	)	,
(	574	)	,
(	576	)	,
(	578	)	,
(	580	)	,
(	583	)	,
(	585	)	,
(	587	)	,
(	589	)	,
(	592	)	,
(	594	)	,
(	596	)	,
(	598	)	,
(	601	)	,
(	603	)	,
(	605	)	,
(	608	)	,
(	610	)	,
(	612	)	,
(	615	)	,
(	617	)	,
(	619	)	,
(	622	)	,
(	624	)	,
(	627	)	,
(	629	)	,
(	631	)	,
(	634	)	,
(	636	)	,
(	639	)	,
(	641	)	,
(	644	)	,
(	646	)	,
(	649	)	,
(	651	)	,
(	654	)	,
(	656	)	,
(	659	)	,
(	661	)	,
(	664	)	,
(	667	)	,
(	669	)	,
(	672	)	,
(	674	)	,
(	677	)	,
(	680	)	,
(	682	)	,
(	685	)	,
(	688	)	,
(	690	)	,
(	693	)	,
(	696	)	,
(	698	)	,
(	701	)	,
(	704	)	,
(	706	)	,
(	709	)	,
(	712	)	,
(	715	)	,
(	717	)	,
(	720	)	,
(	723	)	,
(	726	)	,
(	729	)	,
(	731	)	,
(	734	)	,
(	737	)	,
(	740	)	,
(	743	)	,
(	746	)	,
(	749	)	,
(	752	)	,
(	755	)	,
(	757	)	,
(	760	)	,
(	763	)	,
(	766	)	,
(	769	)	,
(	772	)	,
(	775	)	,
(	778	)	,
(	781	)	,
(	784	)	,
(	787	)	,
(	790	)	,
(	793	)	,
(	797	)	,
(	800	)	,
(	803	)	,
(	806	)	,
(	809	)	,
(	812	)	,
(	815	)	,
(	818	)	,
(	822	)	,
(	825	)	,
(	828	)	,
(	831	)	,
(	834	)	,
(	838	)	,
(	841	)	,
(	844	)	,
(	847	)	,
(	851	)	,
(	854	)	,
(	857	)	,
(	860	)	,
(	864	)	,
(	867	)	,
(	870	)	,
(	874	)	,
(	877	)	,
(	880	)	,
(	884	)	,
(	887	)	,
(	891	)	,
(	894	)	,
(	898	)	,
(	901	)	,
(	904	)	,
(	908	)	,
(	911	)	,
(	915	)	,
(	918	)	,
(	922	)	,
(	925	)	,
(	929	)	,
(	933	)	,
(	936	)	,
(	940	)	,
(	943	)	,
(	947	)	,
(	951	)	,
(	954	)	,
(	958	)	,
(	961	)	,
(	965	)	,
(	969	)	,
(	973	)	,
(	976	)	,
(	980	)	,
(	984	)	,
(	987	)	,
(	991	)	,
(	995	)	,
(	999	)	,
(	1002	)	,
(	1006	)	,
(	1010	)	,
(	1014	)	,
(	1018	)	,
(	1022	)	,
(	1026	)	,
(	1029	)	,
(	1033	)	,
(	1037	)	,
(	1041	)	,
(	1045	)	,
(	1049	)	,
(	1053	)	,
(	1057	)	,
(	1061	)	,
(	1065	)	,
(	1069	)	,
(	1073	)	,
(	1077	)	,
(	1081	)	,
(	1085	)	,
(	1089	)	,
(	1093	)	,
(	1097	)	,
(	1101	)	,
(	1106	)	,
(	1110	)	,
(	1114	)	,
(	1118	)	,
(	1122	)	,
(	1126	)	,
(	1131	)	,
(	1135	)	,
(	1139	)	,
(	1143	)	,
(	1148	)	,
(	1152	)	,
(	1156	)	,
(	1160	)	,
(	1165	)	,
(	1169	)	,
(	1173	)	,
(	1178	)	,
(	1182	)	,
(	1187	)	,
(	1191	)	,
(	1195	)	,
(	1200	)	,
(	1204	)	,
(	1209	)	,
(	1213	)	,
(	1218	)	,
(	1222	)	,
(	1227	)	,
(	1231	)	,
(	1236	)	,
(	1240	)	,
(	1245	)	,
(	1249	)	,
(	1254	)	,
(	1259	)	,
(	1263	)	,
(	1268	)	,
(	1272	)	,
(	1277	)	,
(	1282	)	,
(	1287	)	,
(	1291	)	,
(	1296	)	,
(	1301	)	,
(	1305	)	,
(	1310	)	,
(	1315	)	,
(	1320	)	,
(	1325	)	,
(	1329	)	,
(	1334	)	,
(	1339	)	,
(	1344	)	,
(	1349	)	,
(	1354	)	,
(	1359	)	,
(	1363	)	,
(	1368	)	,
(	1373	)	,
(	1378	)	,
(	1383	)	,
(	1388	)	,
(	1393	)	,
(	1398	)	,
(	1403	)	,
(	1408	)	,
(	1413	)	,
(	1419	)	,
(	1424	)	,
(	1429	)	,
(	1434	)	,
(	1439	)	,
(	1444	)	,
(	1449	)	,
(	1455	)	,
(	1460	)	,
(	1465	)	,
(	1470	)	,
(	1475	)	,
(	1481	)	,
(	1486	)	,
(	1491	)	,
(	1497	)	,
(	1502	)	,
(	1507	)	,
(	1513	)	,
(	1518	)	,
(	1523	)	,
(	1529	)	,
(	1534	)	,
(	1539	)	,
(	1545	)	,
(	1550	)	,
(	1556	)	,
(	1561	)	,
(	1567	)	,
(	1572	)	,
(	1578	)	,
(	1583	)	,
(	1589	)	,
(	1595	)	,
(	1600	)	,
(	1606	)	,
(	1611	)	,
(	1617	)	,
(	1623	)	,
(	1628	)	,
(	1634	)	,
(	1640	)	,
(	1645	)	,
(	1651	)	,
(	1657	)	,
(	1663	)	,
(	1669	)	,
(	1674	)	,
(	1680	)	,
(	1686	)	,
(	1692	)	,
(	1698	)	,
(	1704	)	,
(	1709	)	,
(	1715	)	,
(	1721	)	,
(	1727	)	,
(	1733	)	,
(	1739	)	,
(	1745	)	,
(	1751	)	,
(	1757	)	,
(	1763	)	,
(	1769	)	,
(	1775	)	,
(	1781	)	,
(	1788	)	,
(	1794	)	,
(	1800	)	,
(	1806	)	,
(	1812	)	,
(	1818	)	,
(	1825	)	,
(	1831	)	,
(	1837	)	,
(	1843	)	,
(	1850	)	,
(	1856	)	,
(	1862	)	,
(	1868	)	,
(	1875	)	,
(	1881	)	,
(	1887	)	,
(	1894	)	,
(	1900	)	,
(	1907	)	,
(	1913	)	,
(	1920	)	,
(	1926	)	,
(	1933	)	,
(	1939	)	,
(	1946	)	,
(	1952	)	,
(	1959	)	,
(	1965	)	,
(	1972	)	,
(	1978	)	,
(	1985	)	,
(	1992	)	,
(	1998	)	,
(	2005	)	,
(	2012	)	,
(	2018	)	,
(	2025	)	,
(	2032	)	,
(	2039	)	,
(	2045	)	,
(	2052	)	,
(	2059	)	,
(	2066	)	,
(	2073	)	,
(	2080	)	,
(	2086	)	,
(	2093	)	,
(	2100	)	,
(	2107	)	,
(	2114	)	,
(	2121	)	,
(	2128	)	,
(	2135	)	,
(	2142	)	,
(	2149	)	,
(	2156	)	,
(	2163	)	,
(	2170	)	,
(	2178	)	,
(	2185	)	,
(	2192	)	,
(	2199	)	,
(	2206	)	,
(	2213	)	,
(	2221	)	,
(	2228	)	,
(	2235	)	,
(	2242	)	,
(	2250	)	,
(	2257	)	,
(	2264	)	,
(	2272	)	,
(	2279	)	,
(	2286	)	,
(	2294	)	,
(	2301	)	,
(	2309	)	,
(	2316	)	,
(	2324	)	,
(	2331	)	,
(	2339	)	,
(	2346	)	,
(	2354	)	,
(	2361	)	,
(	2369	)	,
(	2376	)	,
(	2384	)	,
(	2392	)	,
(	2399	)	,
(	2407	)	,
(	2415	)	,
(	2422	)	,
(	2430	)	,
(	2438	)	,
(	2446	)	,
(	2454	)	,
(	2461	)	,
(	2469	)	,
(	2477	)	,
(	2485	)	,
(	2493	)	,
(	2501	)	,
(	2509	)	,
(	2517	)	,
(	2525	)	,
(	2532	)	,
(	2540	)	,
(	2549	)	,
(	2557	)	,
(	2565	)	,
(	2573	)	,
(	2581	)	,
(	2589	)	,
(	2597	)	,
(	2605	)	,
(	2613	)	,
(	2622	)	,
(	2630	)	,
(	2638	)	,
(	2646	)	,
(	2655	)	,
(	2663	)	,
(	2671	)	,
(	2679	)	,
(	2688	)	,
(	2696	)	,
(	2705	)	,
(	2713	)	,
(	2721	)	,
(	2730	)	,
(	2738	)	,
(	2747	)	,
(	2755	)	,
(	2764	)	,
(	2772	)	,
(	2781	)	,
(	2789	)	,
(	2798	)	,
(	2807	)	,
(	2815	)	,
(	2824	)	,
(	2833	)	,
(	2841	)	,
(	2850	)	,
(	2859	)	,
(	2868	)	,
(	2876	)	,
(	2885	)	,
(	2894	)	,
(	2903	)	,
(	2912	)	,
(	2921	)	,
(	2930	)	,
(	2938	)	,
(	2947	)	,
(	2956	)	,
(	2965	)	,
(	2974	)	,
(	2983	)	,
(	2992	)	,
(	3002	)	,
(	3011	)	,
(	3020	)	,
(	3029	)	,
(	3038	)	,
(	3047	)	,
(	3056	)	,
(	3066	)	,
(	3075	)	,
(	3084	)	,
(	3093	)	,
(	3103	)	,
(	3112	)	,
(	3121	)	,
(	3131	)	,
(	3140	)	,
(	3149	)	,
(	3159	)	,
(	3168	)	,
(	3178	)	,
(	3187	)	,
(	3197	)	,
(	3206	)	,
(	3216	)	,
(	3225	)	,
(	3235	)	,
(	3245	)	,
(	3254	)	,
(	3264	)	,
(	3274	)	,
(	3283	)	,
(	3293	)	,
(	3303	)	,
(	3313	)	,
(	3322	)	,
(	3332	)	,
(	3342	)	,
(	3352	)	,
(	3362	)	,
(	3372	)	,
(	3381	)	,
(	3391	)	,
(	3401	)	,
(	3411	)	,
(	3421	)	,
(	3431	)	,
(	3441	)	,
(	3451	)	,
(	3462	)	,
(	3472	)	,
(	3482	)	,
(	3492	)	,
(	3502	)	,
(	3512	)	,
(	3523	)	,
(	3533	)	,
(	3543	)	,
(	3553	)	,
(	3564	)	,
(	3574	)	,
(	3584	)	,
(	3595	)	,
(	3605	)	,
(	3616	)	,
(	3626	)	,
(	3636	)	,
(	3647	)	,
(	3657	)	,
(	3668	)	,
(	3678	)	,
(	3689	)	,
(	3700	)	,
(	3710	)	,
(	3721	)	,
(	3732	)	,
(	3742	)	,
(	3753	)	,
(	3764	)	,
(	3774	)	,
(	3785	)	,
(	3796	)	,
(	3807	)	,
(	3818	)	,
(	3829	)	,
(	3840	)	,
(	3850	)	,
(	3861	)	,
(	3872	)	,
(	3883	)	,
(	3894	)	,
(	3905	)	,
(	3916	)	,
(	3927	)	,
(	3939	)	,
(	3950	)	,
(	3961	)	,
(	3972	)	,
(	3983	)	,
(	3994	)	,
(	4006	)	,
(	4017	)	,
(	4028	)	,
(	4040	)	,
(	4051	)	,
(	4062	)	,
(	4074	)	,
(	4085	)	,
(	4096	)	,
(	4108	)	,
(	4119	)	,
(	4131	)	,
(	4142	)	,
(	4154	)	,
(	4166	)	,
(	4177	)	,
(	4189	)	,
(	4200	)	,
(	4212	)	,
(	4224	)	,
(	4235	)	,
(	4247	)	,
(	4259	)	,
(	4271	)	,
(	4283	)	,
(	4294	)	,
(	4306	)	,
(	4318	)	,
(	4330	)	,
(	4342	)	,
(	4354	)	,
(	4366	)	,
(	4378	)	,
(	4390	)	,
(	4402	)	,
(	4414	)	,
(	4426	)	,
(	4438	)	,
(	4450	)	,
(	4463	)	,
(	4475	)	,
(	4487	)	,
(	4499	)	,
(	4512	)	,
(	4524	)	,
(	4536	)	,
(	4548	)	,
(	4561	)	,
(	4573	)	,
(	4586	)	,
(	4598	)	,
(	4611	)	,
(	4623	)	,
(	4636	)	,
(	4648	)	,
(	4661	)	,
(	4673	)	,
(	4686	)	,
(	4699	)	,
(	4711	)	,
(	4724	)	,
(	4737	)	,
(	4749	)	,
(	4762	)	,
(	4775	)	,
(	4788	)	,
(	4801	)	,
(	4814	)	,
(	4826	)	,
(	4839	)	,
(	4852	)	,
(	4865	)	,
(	4878	)	,
(	4891	)	,
(	4904	)	,
(	4917	)	,
(	4931	)	,
(	4944	)	,
(	4957	)	,
(	4970	)	,
(	4983	)	,
(	4996	)	,
(	5010	)	,
(	5023	)	,
(	5036	)	,
(	5050	)	,
(	5063	)	,
(	5076	)	,
(	5090	)	,
(	5103	)	,
(	5117	)	,
(	5130	)	,
(	5144	)	,
(	5157	)	,
(	5171	)	,
(	5184	)	,
(	5198	)	,
(	5212	)	,
(	5225	)	,
(	5239	)	,
(	5253	)	,
(	5266	)	,
(	5280	)	,
(	5294	)	,
(	5308	)	,
(	5322	)	,
(	5336	)	,
(	5350	)	,
(	5363	)	,
(	5377	)	,
(	5391	)	,
(	5405	)	,
(	5419	)	,
(	5434	)	,
(	5448	)	,
(	5462	)	,
(	5476	)	,
(	5490	)	,
(	5504	)	,
(	5519	)	,
(	5533	)	,
(	5547	)	,
(	5561	)	,
(	5576	)	,
(	5590	)	,
(	5604	)	,
(	5619	)	,
(	5633	)	,
(	5648	)	,
(	5662	)	,
(	5677	)	,
(	5691	)	,
(	5706	)	,
(	5721	)	,
(	5735	)	,
(	5750	)	,
(	5765	)	,
(	5779	)	,
(	5794	)	,
(	5809	)	,
(	5824	)	,
(	5838	)	,
(	5853	)	,
(	5868	)	,
(	5883	)	,
(	5898	)	,
(	5913	)	,
(	5928	)	,
(	5943	)	,
(	5958	)	,
(	5973	)	,
(	5988	)	,
(	6003	)	,
(	6019	)	,
(	6034	)	,
(	6049	)	,
(	6064	)	,
(	6080	)	,
(	6095	)	,
(	6110	)	,
(	6126	)	,
(	6141	)	,
(	6156	)	,
(	6172	)	,
(	6187	)	,
(	6203	)	,
(	6218	)	,
(	6234	)	,
(	6250	)	,
(	6265	)	,
(	6281	)	,
(	6296	)	,
(	6312	)	,
(	6328	)	,
(	6344	)	,
(	6359	)	,
(	6375	)	,
(	6391	)	,
(	6407	)	,
(	6423	)	,
(	6439	)	,
(	6455	)	,
(	6471	)	,
(	6487	)	,
(	6503	)	,
(	6519	)	,
(	6535	)	,
(	6551	)	,
(	6567	)	,
(	6584	)	,
(	6600	)	,
(	6616	)	,
(	6632	)	,
(	6649	)	,
(	6665	)	,
(	6681	)	,
(	6698	)	,
(	6714	)	,
(	6731	)	,
(	6747	)	,
(	6764	)	,
(	6780	)	,
(	6797	)	,
(	6813	)	,
(	6830	)	,
(	6847	)	,
(	6863	)	,
(	6880	)	,
(	6897	)	,
(	6914	)	,
(	6930	)	,
(	6947	)	,
(	6964	)	,
(	6981	)	,
(	6998	)	,
(	7015	)	,
(	7032	)	,
(	7049	)	,
(	7066	)	,
(	7083	)	,
(	7100	)	,
(	7117	)	,
(	7135	)	,
(	7152	)	,
(	7169	)	,
(	7186	)	,
(	7204	)	,
(	7221	)	,
(	7238	)	,
(	7256	)	,
(	7273	)	,
(	7291	)	,
(	7308	)	,
(	7326	)	,
(	7343	)	,
(	7361	)	,
(	7378	)	,
(	7396	)	,
(	7414	)	,
(	7431	)	,
(	7449	)	,
(	7467	)	,
(	7484	)	,
(	7502	)	,
(	7520	)	,
(	7538	)	,
(	7556	)	,
(	7574	)	,
(	7592	)	,
(	7610	)	,
(	7628	)	,
(	7646	)	,
(	7664	)	,
(	7682	)	,
(	7700	)	,
(	7719	)	,
(	7737	)	,
(	7755	)	,
(	7773	)	,
(	7792	)	,
(	7810	)	,
(	7828	)	,
(	7847	)	,
(	7865	)	,
(	7884	)	,
(	7902	)	,
(	7921	)	,
(	7939	)	,
(	7958	)	,
(	7977	)	,
(	7995	)	,
(	8014	)	,
(	8033	)	,
(	8051	)	,
(	8070	)	,
(	8089	)	,
(	8108	)	,
(	8127	)	,
(	8146	)	,
(	8165	)	,
(	8184	)	,
(	8203	)	,
(	8222	)	,
(	8241	)	,
(	8260	)	,
(	8279	)	,
(	8298	)	,
(	8318	)	,
(	8337	)	,
(	8356	)	,
(	8375	)	,
(	8395	)	,
(	8414	)	,
(	8433	)	,
(	8453	)	,
(	8472	)	,
(	8492	)	,
(	8511	)	,
(	8531	)	,
(	8551	)	,
(	8570	)	,
(	8590	)	,
(	8610	)	,
(	8629	)	,
(	8649	)	,
(	8669	)	,
(	8689	)	,
(	8709	)	,
(	8729	)	,
(	8748	)	,
(	8768	)	,
(	8788	)	,
(	8809	)	,
(	8829	)	,
(	8849	)	,
(	8869	)	,
(	8889	)	,
(	8909	)	,
(	8929	)	,
(	8950	)	,
(	8970	)	,
(	8990	)	,
(	9011	)	,
(	9031	)	,
(	9052	)	,
(	9072	)	,
(	9093	)	,
(	9113	)	,
(	9134	)	,
(	9154	)	,
(	9175	)	,
(	9196	)	,
(	9216	)	,
(	9237	)	,
(	9258	)	,
(	9279	)	,
(	9299	)	,
(	9320	)	,
(	9341	)	,
(	9362	)	,
(	9383	)	,
(	9404	)	,
(	9425	)	,
(	9446	)	,
(	9467	)	,
(	9489	)	,
(	9510	)	,
(	9531	)	,
(	9552	)	,
(	9574	)	,
(	9595	)	,
(	9616	)	,
(	9638	)	,
(	9659	)	,
(	9681	)	,
(	9702	)	,
(	9724	)	,
(	9745	)	,
(	9767	)	,
(	9788	)	,
(	9810	)	,
(	9832	)	,
(	9854	)	,
(	9875	)	,
(	9897	)	,
(	9919	)	,
(	9941	)	,
(	9963	)	,
(	9985	)	,
(	10007	)	,
(	10029	)	,
(	10051	)	,
(	10073	)	,
(	10095	)	,
(	10117	)	,
(	10139	)	,
(	10162	)	,
(	10184	)	,
(	10206	)	,
(	10229	)	,
(	10251	)	,
(	10273	)	,
(	10296	)	,
(	10318	)	,
(	10341	)	,
(	10363	)	,
(	10386	)	,
(	10409	)	,
(	10431	)	,
(	10454	)	,
(	10477	)	,
(	10500	)	,
(	10522	)	,
(	10545	)	,
(	10568	)	,
(	10591	)	,
(	10614	)	,
(	10637	)	,
(	10660	)	,
(	10683	)	,
(	10706	)	,
(	10729	)	,
(	10753	)	,
(	10776	)	,
(	10799	)	,
(	10822	)	,
(	10846	)	,
(	10869	)	,
(	10892	)	,
(	10916	)	,
(	10939	)	,
(	10963	)	,
(	10986	)	,
(	11010	)	,
(	11034	)	,
(	11057	)	,
(	11081	)	,
(	11105	)	,
(	11128	)	,
(	11152	)	,
(	11176	)	,
(	11200	)	,
(	11224	)	,
(	11248	)	,
(	11272	)	,
(	11296	)	,
(	11320	)	,
(	11344	)	,
(	11368	)	,
(	11392	)	,
(	11416	)	,
(	11441	)	,
(	11465	)	,
(	11489	)	,
(	11514	)	,
(	11538	)	,
(	11563	)	,
(	11587	)	,
(	11612	)	,
(	11636	)	,
(	11661	)	,
(	11685	)	,
(	11710	)	,
(	11735	)	,
(	11759	)	,
(	11784	)	,
(	11809	)	,
(	11834	)	,
(	11859	)	,
(	11884	)	,
(	11909	)	,
(	11934	)	,
(	11959	)	,
(	11984	)	,
(	12009	)	,
(	12034	)	,
(	12059	)	,
(	12085	)	,
(	12110	)	,
(	12135	)	,
(	12160	)	,
(	12186	)	,
(	12211	)	,
(	12237	)	,
(	12262	)	,
(	12288	)	,
(	12313	)	,
(	12339	)	,
(	12365	)	,
(	12390	)	,
(	12416	)	,
(	12442	)	,
(	12468	)	,
(	12494	)	,
(	12520	)	,
(	12545	)	,
(	12571	)	,
(	12597	)	,
(	12624	)	,
(	12650	)	,
(	12676	)	,
(	12702	)	,
(	12728	)	,
(	12754	)	,
(	12781	)	,
(	12807	)	,
(	12833	)	,
(	12860	)	,
(	12886	)	,
(	12913	)	,
(	12939	)	,
(	12966	)	,
(	12993	)	,
(	13019	)	,
(	13046	)	,
(	13073	)	,
(	13099	)	,
(	13126	)	,
(	13153	)	,
(	13180	)	,
(	13207	)	,
(	13234	)	,
(	13261	)	,
(	13288	)	,
(	13315	)	,
(	13342	)	,
(	13369	)	,
(	13396	)	,
(	13424	)	,
(	13451	)	,
(	13478	)	,
(	13506	)	,
(	13533	)	,
(	13561	)	,
(	13588	)	,
(	13616	)	,
(	13643	)	,
(	13671	)	,
(	13699	)	,
(	13726	)	,
(	13754	)	,
(	13782	)	,
(	13810	)	,
(	13837	)	,
(	13865	)	,
(	13893	)	,
(	13921	)	,
(	13949	)	,
(	13977	)	,
(	14005	)	,
(	14034	)	,
(	14062	)	,
(	14090	)	,
(	14118	)	,
(	14147	)	,
(	14175	)	,
(	14203	)	,
(	14232	)	,
(	14260	)	,
(	14289	)	,
(	14317	)	,
(	14346	)	,
(	14375	)	,
(	14403	)	,
(	14432	)	,
(	14461	)	,
(	14490	)	,
(	14519	)	,
(	14547	)	,
(	14576	)	,
(	14605	)	,
(	14634	)	,
(	14664	)	,
(	14693	)	,
(	14722	)	,
(	14751	)	,
(	14780	)	,
(	14809	)	,
(	14839	)	,
(	14868	)	,
(	14898	)	,
(	14927	)	,
(	14957	)	,
(	14986	)	,
(	15016	)	,
(	15045	)	,
(	15075	)	,
(	15105	)	,
(	15134	)	,
(	15164	)	,
(	15194	)	,
(	15224	)	,
(	15254	)	,
(	15284	)	,
(	15314	)	,
(	15344	)	,
(	15374	)	,
(	15404	)	,
(	15434	)	,
(	15464	)	,
(	15495	)	,
(	15525	)	,
(	15555	)	,
(	15586	)	,
(	15616	)	,
(	15647	)	,
(	15677	)	,
(	15708	)	,
(	15738	)	,
(	15769	)	,
(	15800	)	,
(	15831	)	,
(	15861	)	,
(	15892	)	,
(	15923	)	,
(	15954	)	,
(	15985	)	,
(	16016	)	,
(	16047	)	,
(	16078	)	,
(	16109	)	,
(	16140	)	,
(	16172	)	,
(	16203	)	,
(	16234	)	,
(	16266	)	,
(	16297	)	,
(	16328	)	,
(	16360	)	,
(	16391	)	,
(	16423	)	,
(	16455	)	,
(	16486	)	,
(	16518	)	,
(	16550	)	,
(	16582	)	,
(	16613	)	,
(	16645	)	,
(	16677	)	,
(	16709	)	,
(	16741	)	,
(	16773	)	,
(	16805	)	,
(	16838	)	,
(	16870	)	,
(	16902	)	,
(	16934	)	,
(	16967	)	,
(	16999	)	,
(	17032	)	,
(	17064	)	,
(	17097	)	




);


end package LUT_pkg;
